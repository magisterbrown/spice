inverter circuit
.model nmfeet nmos ()
.model pmfeet pmos ()

Vcc cc 0 2
V1 ain 0 pulse (0 2 5n 2n 2n 90n 180n)
V2 bin 0 pulse (0 2 5n 2n 2n 45n 80n)

Mnmos1 nm1out ain 0 0 nmfeet
Mnmos2 out bin nm1out 0 nmfeet

Mpmos1 out ain cc cc pmfeet
Mpmos2 out bin cc cc pmfeet


.control
    tran 100p 150n
    print out ain bin
    exit
.endc
.end
